module LZC (
  input
  output
);

endmodule
